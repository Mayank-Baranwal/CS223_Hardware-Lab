`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:49:45 02/08/2019 
// Design Name: 
// Module Name:    CLA_16bit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module CLA_16bit(
    input [15:0] A,B,
	 input Cin,
	 output [15:0] C,S,
	 output Cout
	 );

	wire G0,G4,G8,G12;
	wire P0,P4,P8,P12;
	
endmodule
